package `VITISNETP4_VERIF_PKG_NAME;

   `include `"`VITISNETP4_AGENT_INCLUDE_FILE`"

endpackage : `VITISNETP4_VERIF_PKG_NAME

