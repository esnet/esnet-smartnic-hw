package p4_and_verilog_pkg;
    // --------------------------------------------------------------
    // Imports
    // --------------------------------------------------------------
    import sdnet_0_pkg::*;

    // --------------------------------------------------------------
    // Parameters & Typedefs
    // --------------------------------------------------------------
    // User metadata
    typedef USER_META_DATA_T user_metadata_t;

endpackage : p4_and_verilog_pkg
