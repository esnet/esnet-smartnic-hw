package smartnic_322mhz_app_pkg;

    localparam bit INCLUDE_HBM = 1'b1;

endpackage : smartnic_322mhz_app_pkg
