package xilinx_alveo_au250_pkg;

    // --------------------------------------------------------------
    // Parameters
    // --------------------------------------------------------------
    localparam int PCIE_LINK_WID = 16;
    localparam int NUM_QSFP = 2;

endpackage : xilinx_alveo_au250_pkg
