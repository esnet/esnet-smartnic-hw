../../../../../../src/vitisnetp4/verif/src/vitisnetp4_verif_pkg.sv