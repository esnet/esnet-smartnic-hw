package tb_pkg;
    import axi4l_verif_pkg::*;
    import axi4s_verif_pkg::*;
    import p4_app_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "timestamp_agent.svh"
    `include "tb_env.svh"

endpackage : tb_pkg
