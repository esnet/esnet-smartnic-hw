package smartnic_verif_pkg;

   `include "smartnic_model.svh"

endpackage : smartnic_verif_pkg
