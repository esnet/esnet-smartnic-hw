`include "svunit_defines.svh"

//===================================
// (Failsafe) timeout
//===================================
`define SVUNIT_TIMEOUT 200us

module smartnic_322mhz_datapath_unit_test;

    // Testcase name
    string name = "smartnic_322mhz_datapath_ut";

    // SVUnit base testcase
    svunit_pkg::svunit_testcase svunit_ut;

    //===================================
    // DUT + testbench
    //===================================
    // This test suite references the common smartnic_322mhz
    // testbench top level. The 'tb' module is
    // loaded into the tb_glbl scope, so is available
    // at tb_glbl.tb.
    //
    // Interaction with the testbench is expected to occur
    // via the testbench environment class (tb_env). A
    // reference to the testbench environment is provided
    // here for convenience.
    tb_pkg::tb_env env;

    //===================================
    // Import common testcase tasks
    //=================================== 
    `include "../../tests/common/tasks.svh"
       
    //===================================
    // Connect AXI-S sample interface
    //===================================

    /*
    assign tb.axis_sample_clk = tb.clk;
    assign tb.axis_sample_aresetn = !tb.rst;
    assign tb.axis_sample_if.tvalid = tb.DUT.bypass_mux_to_switch.axi4s_in.tvalid;
    assign tb.axis_sample_if.tlast  = tb.DUT.bypass_mux_to_switch.axi4s_in.tlast;
    assign tb.axis_sample_if.tdata  = tb.DUT.bypass_mux_to_switch.axi4s_in.tdata;
    assign tb.axis_sample_if.tkeep  = tb.DUT.bypass_mux_to_switch.axi4s_in.tkeep;
    assign tb.axis_sample_if.tuser  = tb.DUT.bypass_mux_to_switch.axi4s_in.tuser;
    assign tb.axis_sample_if.tready = tb.DUT.bypass_mux_to_switch.axi4s_in.tready;
    */

    //===================================
    // Build
    //===================================
    function void build();
        svunit_ut = new(name);

        // Build testbench
        tb.build();

        // Retrieve reference to testbench environment class
        env = tb.env;

    endfunction

    //===================================
    // Global test variables
    //===================================
    localparam NUM_PORTS = 4;
    localparam FIFO_DEPTH = 410.0; // 124 (fifo_async) + 2 x 143 (axi4s_pkt_discard_ovfl)

    smartnic_322mhz_reg_pkg::reg_port_config_t set_config;

    // variables for switch tests.
    import smartnic_322mhz_pkg::*;
    port_t out_port_map [NUM_PORTS-1:0];  // vector specifies output port for each input stream.

    string in_pcap  [NUM_PORTS-1:0];  // vector specifies the in_pcap file for each input stream.
    string out_pcap [NUM_PORTS-1:0];  // vector specifies the out_pcap file for each input stream.

    // variables for probe checks.
    int tx_pkt_cnt  [NUM_PORTS-1:0];  // captures the tx pkt & byte counts from the pcap file for a given test.
    int tx_byte_cnt [NUM_PORTS-1:0];

    int rx_pkt_cnt  [NUM_PORTS-1:0];  // captures the rx pkt & byte counts from the pcap file for a given test.
    int rx_byte_cnt [NUM_PORTS-1:0];

    int rx_pkt_tot  = 0;
    int rx_byte_tot = 0;

    // variables for discard tests.
    int	pkt_len     [NUM_PORTS-1:0];
    int exp_pkt_cnt [NUM_PORTS-1:0];  // vector specifies the expected number of pkts received for each stream.

   
    //===================================
    // Setup for running the Unit Tests
    //===================================
    task setup();
        // default variable configuration
         in_pcap[0] = "../../../tests/common/pcap/20xrandom_pkts.pcap";
        out_pcap[0] = "../../../tests/common/pcap/20xrandom_pkts.pcap";
         in_pcap[1] = "../../../tests/common/pcap/30xrandom_pkts.pcap";
        out_pcap[1] = "../../../tests/common/pcap/30xrandom_pkts.pcap";
         in_pcap[2] = "../../../tests/common/pcap/40xrandom_pkts.pcap";
        out_pcap[2] = "../../../tests/common/pcap/40xrandom_pkts.pcap";
         in_pcap[3] = "../../../tests/common/pcap/50xrandom_pkts.pcap";
        out_pcap[3] = "../../../tests/common/pcap/50xrandom_pkts.pcap";

        out_port_map = {2'h0, 2'h2, 2'h3, 2'h1};
        pkt_len      = {0, 0, 0, 0};  
        exp_pkt_cnt  = {0, 0, 0, 0};  // if exp_pkt_cnt field is set 0, value is determined from pcap file.

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(0);

        svunit_ut.setup();

        // Issue reset (both datapath and management domains)
        reset();

       // Write port_config register to enable app bypass mode.
        set_config.input_enable  = smartnic_322mhz_reg_pkg::PORT_CONFIG_INPUT_ENABLE_BOTH;
        set_config.output_enable = smartnic_322mhz_reg_pkg::PORT_CONFIG_OUTPUT_ENABLE_USE_META;
        set_config.app_bypass = 1'b1;
        set_config.app_tpause = 1'b0;
        env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);

        `INFO("Waiting to initialize axis fifos...");
        for (integer i = 0; i < 100 ; i=i+1 ) begin
          @(posedge tb.clk);
        end

    endtask


    //===================================
    // Here we deconstruct anything we
    // need after running the Unit Tests
    //===================================
    task teardown();
        `INFO("Waiting to end testcase...");
        for (integer i = 0; i < 100 ; i=i+1 ) @(posedge tb.clk);
        `INFO("Ending testcase!");

        svunit_ut.teardown();

    endtask

    //=======================================================================
    // TESTS
    //=======================================================================

    //===================================
    // All tests are defined between the
    // SVUNIT_TESTS_BEGIN/END macros
    //
    // Each individual test must be
    // defined between `SVTEST(_NAME_)
    // `SVTEST_END
    //
    // i.e.
    //   `SVTEST(mytest)
    //     <test code>
    //   `SVTEST_END
    //===================================

    `SVUNIT_TESTS_BEGIN

    `SVTEST(switch_basic_sanity)
        out_port_map = {2'h3, 2'h2, 2'h1, 2'h0}; 

        run_stream_test(); check_stream_test_probes;
    `SVTEST_END


    `SVTEST(switch_with_halt_probe_counters)
        out_port_map = {2'h1, 2'h2, 2'h0, 2'h3};

        halt_probe_counters;

        run_stream_test();

        check_stream_probes ( .in_port(0), .out_port(out_port_map[0]), .exp_good_pkts(0), .exp_good_bytes(0) );
        check_stream_probes ( .in_port(1), .out_port(out_port_map[1]), .exp_good_pkts(0), .exp_good_bytes(0) );
        check_stream_probes ( .in_port(3), .out_port(out_port_map[3]), .exp_good_pkts(0), .exp_good_bytes(0) );
        check_stream_probes ( .in_port(2), .out_port(out_port_map[2]), .exp_good_pkts(0), .exp_good_bytes(0) );
   
        check_probe ( .base_addr('ha000), .exp_pkt_cnt(0), .exp_byte_cnt(0) );
        check_probe ( .base_addr('ha800), .exp_pkt_cnt(0), .exp_byte_cnt(0) );
    `SVTEST_END


    `SVTEST(switch_with_discards)
         in_pcap[0] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
        out_pcap[0] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
         pkt_len[0] = 1518;
         in_pcap[1] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
        out_pcap[1] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
         pkt_len[1] = 9100;
         in_pcap[2] = "../../../tests/common/pcap/50xrandom_pkts.pcap";
        out_pcap[2] = "../../../tests/common/pcap/50xrandom_pkts.pcap";
         pkt_len[2] = 0;
         in_pcap[3] = "../../../tests/common/pcap/128x566B_pkts.pcap";
        out_pcap[3] = "../../../tests/common/pcap/128x566B_pkts.pcap";
         pkt_len[3] = 566;

        // FIFO holds FIFO_DEPTH x 64B good packets (all others dropped).
        for (int i=0; i<NUM_PORTS; i++)
           exp_pkt_cnt[i] = (pkt_len[i]==0) ? 0 : $ceil(FIFO_DEPTH/$ceil(pkt_len[i]/64.0));

        force tb.axis_out_if[0].tready = 0;  // force backpressure on egress ports with discard points
        force tb.axis_out_if[1].tready = 0;
        force tb.axis_out_if[2].tready = 0;
        force tb.axis_out_if[3].tready = 0;

        env.axis_driver[0].set_min_gap(2*$ceil(pkt_len[0]/64.0));  // set gap to 2 pkts.
        env.axis_driver[1].set_min_gap(2*$ceil(pkt_len[1]/64.0));
        env.axis_driver[2].set_min_gap(2*$ceil(pkt_len[2]/64.0));
        env.axis_driver[3].set_min_gap(2*$ceil(pkt_len[3]/64.0));

        fork
           run_stream_test();

           begin
              #(50us);
              force   tb.axis_out_if[0].tready = 1; release tb.axis_out_if[0].tready;
              force   tb.axis_out_if[1].tready = 1; release tb.axis_out_if[1].tready;
              force   tb.axis_out_if[2].tready = 1; release tb.axis_out_if[2].tready;
              force   tb.axis_out_if[3].tready = 1; release tb.axis_out_if[3].tready;
           end
	join

         check_stream_test_probes;
    `SVTEST_END


    `SVTEST(max_size_discards)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
        end

        // FIFO holds FIFO_DEPTH x 64B good packets (all others dropped).
        for (int i=0; i<NUM_PORTS; i++) begin
            pkt_len[i] = 1518;
            exp_pkt_cnt[i] = $ceil(FIFO_DEPTH/$ceil(pkt_len[i]/64.0));
        end
        exp_pkt_cnt[2] = 0;  // configures exp_pkt_cnt from pcap file.

        force tb.axis_out_if[0].tready = 0;  // force backpressure on egress ports with discard points
        force tb.axis_out_if[1].tready = 0;
        force tb.axis_out_if[2].tready = 0;
        force tb.axis_out_if[3].tready = 0;

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(2*$ceil(pkt_len[i]/64.0)); // set gap to 2 pkts.

        fork
           run_stream_test();

           begin
              #(50us);
              force   tb.axis_out_if[0].tready = 1; release tb.axis_out_if[0].tready;
              force   tb.axis_out_if[1].tready = 1; release tb.axis_out_if[1].tready;
              force   tb.axis_out_if[2].tready = 1; release tb.axis_out_if[1].tready;
              force   tb.axis_out_if[3].tready = 1; release tb.axis_out_if[3].tready;
           end
	join

        check_stream_test_probes;
    `SVTEST_END

      
    `SVTEST(jumbo_size_discards)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
        end

        // FIFO holds FIFO_DEPTH x 64B good packets (all others dropped).
        for (int i=0; i<NUM_PORTS; i++) begin
            pkt_len[i] = 9100;
            exp_pkt_cnt[i] = $ceil(FIFO_DEPTH/$ceil(pkt_len[i]/64.0));
        end
        exp_pkt_cnt[2] = 0;  // configures exp_pkt_cnt from pcap file.

        force tb.axis_out_if[0].tready = 0;  // force backpressure on egress ports with discard points
        force tb.axis_out_if[1].tready = 0;
        force tb.axis_out_if[2].tready = 0;
        force tb.axis_out_if[3].tready = 0;

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(2*$ceil(pkt_len[i]/64.0)); // set gap to 2 pkts.

        fork
           run_stream_test();

           begin
              #(50us);
              force   tb.axis_out_if[0].tready = 1; release tb.axis_out_if[0].tready;
              force   tb.axis_out_if[1].tready = 1; release tb.axis_out_if[1].tready;
              force   tb.axis_out_if[2].tready = 1; release tb.axis_out_if[1].tready;
              force   tb.axis_out_if[3].tready = 1; release tb.axis_out_if[3].tready;
           end
	join

        check_stream_test_probes;
    `SVTEST_END


    `SVTEST(discards_from_cmac)
         in_pcap[0] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
        out_pcap[0] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
         pkt_len[0] = 9100;
         in_pcap[1] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
        out_pcap[1] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
         pkt_len[1] = 1518;

        // FIFO holds FIFO_DEPTH x 64B good packets (all others dropped).
        for (int i=0; i<NUM_PORTS; i++)
           exp_pkt_cnt[i] = (pkt_len[i]==0) ? 0 : $ceil(FIFO_DEPTH/$ceil(pkt_len[i]/64.0));

        // force backpressure on ingress ports (deasserts tready from app core to ingress switch).
        set_config.app_tpause = 1; env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);
   
        fork
           run_stream_test();

           begin
              #(50us);
              // release backpressure on ingress ports
              set_config.app_tpause = 0; env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);
           end
	join

        check_stream_test_probes (.ingress_ovfl_mode(1));
    `SVTEST_END


    `SVTEST(errored_packets)
         for (int i=0; i<2; i++) begin // 2 iterations

            for (int cmac_port=0; cmac_port<2; cmac_port++) begin // foreach cmac port

               env.axis_driver[cmac_port].set_min_gap(i); // set gap to i cycles.

               // send 10 errored packets i.e. with tuser=1
               send_pcap(.pcap_filename ("../../../tests/common/pcap/64B_multiples_10pkts.pcap"),
                         .id(cmac_port), .dest(cmac_port), .user(1));
               // check error counts
               check_err_probes (.in_port(cmac_port), .exp_err_pkts(10), .exp_err_bytes(3520));

               // send and check unerrored packet stream i.e. with tuser=0 (default)
               run_pkt_stream (.in_port(cmac_port), .out_port(cmac_port),
                               .in_pcap  ("../../../tests/common/pcap/64x1518B_pkts.pcap"),
                               .out_pcap ("../../../tests/common/pcap/64x1518B_pkts.pcap"),
                               .tx_pkt_cnt(tx_pkt_cnt[cmac_port]), .tx_byte_cnt(tx_byte_cnt[cmac_port]),
                               .rx_pkt_cnt(rx_pkt_cnt[cmac_port]), .rx_byte_cnt(rx_byte_cnt[cmac_port]) );

               // check stream probe counts
               check_stream_probes (.in_port(cmac_port), .out_port(cmac_port),
                                    .exp_good_pkts(rx_pkt_cnt[cmac_port]), .exp_good_bytes(rx_byte_cnt[cmac_port]),
                                    .exp_ovfl_pkts(0), .exp_ovfl_bytes(0) );
             end

          end
    `SVTEST_END


    `SVTEST(single_packets)
         env.axis_driver[1].set_min_gap(1000); // set gap to 1000 cycles.

         run_pkt_stream ( .in_port(1), .out_port(1), 
                         .in_pcap  ("../../../tests/common/pcap/64B_multiples_10pkts.pcap"),
                         .out_pcap ("../../../tests/common/pcap/64B_multiples_10pkts.pcap"),
                         .tx_pkt_cnt(tx_pkt_cnt[1]), .tx_byte_cnt(tx_byte_cnt[1]),
                         .rx_pkt_cnt(rx_pkt_cnt[1]), .rx_byte_cnt(rx_byte_cnt[1]) );
    `SVTEST_END


    `SVTEST(port_config_0)
        force tb.axis_in_if[0].tdest = 2'h2; // force axis_in_if[0] to direct all traffic to port 2 (HOST_PORT0). 

        // Write port_config register to direct all traffic to CMAC_PORT0
        set_config.input_enable  = smartnic_322mhz_reg_pkg::PORT_CONFIG_INPUT_ENABLE_PORT0;
        set_config.output_enable = smartnic_322mhz_reg_pkg::PORT_CONFIG_OUTPUT_ENABLE_PORT0;

        env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);

        // Run pkt traffic. Expect rx pkts at CMAC_PORT0, as per port_config setting.
        run_pkt_stream ( .in_port(0), .out_port(0), 
                         .in_pcap ("../../../tests/common/pcap/20xrandom_pkts.pcap"),
                         .out_pcap("../../../tests/common/pcap/20xrandom_pkts.pcap"),
                         .tx_pkt_cnt(tx_pkt_cnt[0]), .tx_byte_cnt(tx_byte_cnt[0]),
                         .rx_pkt_cnt(rx_pkt_cnt[0]), .rx_byte_cnt(rx_byte_cnt[0]) );

         release tb.axis_in_if[0].tdest;
    `SVTEST_END

      
    `SVTEST(port_config_1)
        force tb.axis_in_if[0].tdest = 2'h2; // force axis_in_if[0] to direct all traffic to port 2 (HOST_PORT0). 

        // Write port_config register to direct all traffic to CMAC_PORT1
        set_config.input_enable  = smartnic_322mhz_reg_pkg::PORT_CONFIG_INPUT_ENABLE_PORT0;
        set_config.output_enable = smartnic_322mhz_reg_pkg::PORT_CONFIG_OUTPUT_ENABLE_PORT1;

        env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);

        // Run pkt traffic. Expect rx pkts at CMAC_PORT1, as per port_config setting.
        run_pkt_stream ( .in_port(0), .out_port(1), 
                         .in_pcap ("../../../tests/common/pcap/20xrandom_pkts.pcap"),
                         .out_pcap("../../../tests/common/pcap/20xrandom_pkts.pcap"),
                         .tx_pkt_cnt(tx_pkt_cnt[0]), .tx_byte_cnt(tx_byte_cnt[0]),
                         .rx_pkt_cnt(rx_pkt_cnt[0]), .rx_byte_cnt(rx_byte_cnt[0]) );

         release tb.axis_in_if[0].tdest;
    `SVTEST_END


    `SVTEST(port_config_2)
        force tb.axis_in_if[0].tdest = 2'h2; // force axis_in_if[0] to direct all traffic to port 2 (HOST_PORT0). 

        // Write port_config register to direct all traffic to CMAC_PORT0
        set_config.input_enable  = smartnic_322mhz_reg_pkg::PORT_CONFIG_INPUT_ENABLE_PORT0;
        set_config.output_enable = smartnic_322mhz_reg_pkg::PORT_CONFIG_OUTPUT_ENABLE_C2H;

        env.smartnic_322mhz_reg_blk_agent.write_port_config(set_config);

        // Run pkt traffic. Expect rx pkts at HOST_PORT1, as per port_config setting.
        run_pkt_stream ( .in_port(0), .out_port(3), 
                         .in_pcap ("../../../tests/common/pcap/20xrandom_pkts.pcap"), 
                         .out_pcap("../../../tests/common/pcap/20xrandom_pkts.pcap"), 
                         .tx_pkt_cnt(tx_pkt_cnt[0]), .tx_byte_cnt(tx_byte_cnt[0]),
                         .rx_pkt_cnt(rx_pkt_cnt[0]), .rx_byte_cnt(rx_byte_cnt[0]) );

        release tb.axis_in_if[0].tdest;
    `SVTEST_END


    `SVTEST(min_size_stress)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/512x64B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/512x64B_pkts.pcap";
        end

        run_stream_test(); check_stream_test_probes;
    `SVTEST_END


    `SVTEST(max_size_stress)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/64x1518B_pkts.pcap";
        end

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(2*24);  // set gap to 2 pkts.

        run_stream_test(); check_stream_test_probes;

    `SVTEST_END


    `SVTEST(short_pkt)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/256x54B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/256x54B_pkts.pcap";
        end

        run_stream_test(); check_stream_test_probes;
    `SVTEST_END


    `SVTEST(long_pkt)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/16x9100B_pkts.pcap";
        end

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(2*143);  // set gap to 2 pkts.

        run_stream_test(); check_stream_test_probes;
    `SVTEST_END


    `SVTEST(axi4s_tkeep_stress)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/64B_to_319B_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/64B_to_319B_pkts.pcap";
        end

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(5);  // set gap to 5 cycles.

        run_stream_test(); check_stream_test_probes;
    `SVTEST_END

      
    `SVTEST(random_pkt_size)
        for (int i=0; i<NUM_PORTS; i++) begin
            in_pcap[i] = "../../../tests/common/pcap/100xrandom_pkts.pcap";
           out_pcap[i] = "../../../tests/common/pcap/100xrandom_pkts.pcap";
        end

        for (int i=0; i<NUM_PORTS; i++) env.axis_driver[i].set_min_gap(2*143);  // set gap to 2 jumbo pkts.

        run_stream_test(); check_stream_test_probes;

    `SVTEST_END

    `SVUNIT_TESTS_END



   
    task run_stream_test (input int tpause = 0, twait = 0);
        fork
           run_pkt_stream ( .in_port(0), .out_port(out_port_map[0]), .in_pcap(in_pcap[0]), .out_pcap(out_pcap[0]),
                            .tx_pkt_cnt(tx_pkt_cnt[0]), .tx_byte_cnt(tx_byte_cnt[0]), 
                            .rx_pkt_cnt(rx_pkt_cnt[0]), .rx_byte_cnt(rx_byte_cnt[0]),
                            .exp_pkt_cnt(exp_pkt_cnt[0]),
                            .tpause(tpause), .twait(twait) );

           run_pkt_stream ( .in_port(1), .out_port(out_port_map[1]), .in_pcap(in_pcap[1]), .out_pcap(out_pcap[1]),
                            .tx_pkt_cnt(tx_pkt_cnt[1]), .tx_byte_cnt(tx_byte_cnt[1]), 
                            .rx_pkt_cnt(rx_pkt_cnt[1]), .rx_byte_cnt(rx_byte_cnt[1]),
                            .exp_pkt_cnt(exp_pkt_cnt[1]),
                            .tpause(tpause), .twait(twait) );

           run_pkt_stream ( .in_port(2), .out_port(out_port_map[2]), .in_pcap(in_pcap[2]), .out_pcap(out_pcap[2]),
                            .tx_pkt_cnt(tx_pkt_cnt[2]), .tx_byte_cnt(tx_byte_cnt[2]), 
                            .rx_pkt_cnt(rx_pkt_cnt[2]), .rx_byte_cnt(rx_byte_cnt[2]),
                            .exp_pkt_cnt(exp_pkt_cnt[2]),
                            .tpause(tpause), .twait(twait) );

           run_pkt_stream ( .in_port(3), .out_port(out_port_map[3]), .in_pcap(in_pcap[3]), .out_pcap(out_pcap[3]),
                            .tx_pkt_cnt(tx_pkt_cnt[3]), .tx_byte_cnt(tx_byte_cnt[3]), 
                            .rx_pkt_cnt(rx_pkt_cnt[3]), .rx_byte_cnt(rx_byte_cnt[3]),
                            .exp_pkt_cnt(exp_pkt_cnt[3]),
                            .tpause(tpause), .twait(twait) );

        join
    endtask
   

    task check_stream_test_probes (input logic ingress_ovfl_mode = 0);
        for (int i=0; i<NUM_PORTS; i++) begin
           check_stream_probes (
              .in_port         (i), 
              .out_port        (out_port_map[i]),
              .exp_good_pkts   (rx_pkt_cnt[i]), 
              .exp_good_bytes  (rx_byte_cnt[i]), 
              .exp_ovfl_pkts   (tx_pkt_cnt[i]  - rx_pkt_cnt[i]), 
              .exp_ovfl_bytes  (tx_byte_cnt[i] - rx_byte_cnt[i]),
              .ingress_ovfl_mode   (ingress_ovfl_mode)
           );
	end
    endtask;


    typedef enum logic [31:0] {
        PROBE_FROM_CMAC_PORT0      = 'h8000,
        DROPS_OVFL_FROM_CMAC_PORT0 = 'h8400,
        DROPS_ERR_FROM_CMAC_PORT0  = 'h8800,
        PROBE_FROM_CMAC_PORT1      = 'h8c00,
        DROPS_OVFL_FROM_CMAC_PORT1 = 'h9000,
        DROPS_ERR_FROM_CMAC_PORT1  = 'h9400,
        PROBE_FROM_HOST_PORT0      = 'h9800,
        PROBE_FROM_HOST_PORT1      = 'h9c00,

        PROBE_TO_CMAC_PORT0        = 'hb000,
        DROPS_OVFL_TO_CMAC_PORT0   = 'hb400,
        PROBE_TO_CMAC_PORT1        = 'hb800,
        DROPS_OVFL_TO_CMAC_PORT1   = 'hbc00,
        PROBE_TO_HOST_PORT0        = 'hc000,
        DROPS_OVFL_TO_HOST_PORT0   = 'hc400,
        PROBE_TO_HOST_PORT1        = 'hc800,
        DROPS_OVFL_TO_HOST_PORT1   = 'hcc00
    } cntr_addr_encoding_t;

    typedef union packed {
        cntr_addr_encoding_t  encoded;
        logic [31:0]          raw;
    } cntr_addr_t;

   
    task check_stream_probes ( input port_t       in_port, out_port,
                               input logic [63:0] exp_good_pkts, exp_good_bytes, exp_ovfl_pkts=0, exp_ovfl_bytes=0,
                               input logic        ingress_ovfl_mode = 0 );

        cntr_addr_t in_port_base_addr, out_port_base_addr;
        logic [63:0] exp_tot_pkts, exp_tot_bytes;

        // establish base addr for ingress probe
        case (in_port)
               CMAC_PORT0 : in_port_base_addr = 'h8000;
               CMAC_PORT1 : in_port_base_addr = 'h8c00;
               HOST_PORT0 : in_port_base_addr = 'h9800;
               HOST_PORT1 : in_port_base_addr = 'h9c00;
	    default : in_port_base_addr = 'hxxxx;
        endcase

        // establish base addr for egress probe
        case (out_port)
               CMAC_PORT0 : out_port_base_addr = 'hb000;
               CMAC_PORT1 : out_port_base_addr = 'hb800;
               HOST_PORT0 : out_port_base_addr = 'hc000;
               HOST_PORT1 : out_port_base_addr = 'hc800;
	    default : out_port_base_addr = 'hxxxx;
        endcase

        // establish pkt and byte totals       
        exp_tot_pkts  = exp_good_pkts  + exp_ovfl_pkts;
        exp_tot_bytes = exp_good_bytes + exp_ovfl_bytes;


        // check ingress and egress probe counts
        if (ingress_ovfl_mode)
           check_probe (.base_addr(in_port_base_addr), .exp_pkt_cnt(exp_good_pkts), .exp_byte_cnt(exp_good_bytes));
        else
           check_probe (.base_addr(in_port_base_addr), .exp_pkt_cnt(exp_tot_pkts),  .exp_byte_cnt(exp_tot_bytes));

        check_probe (.base_addr(out_port_base_addr), .exp_pkt_cnt(exp_good_pkts), .exp_byte_cnt(exp_good_bytes));


        // check ingress and egress ovfl counts
        if ( (in_port != HOST_PORT0) && (in_port != HOST_PORT1) ) begin  // no ovfl counters for these ingress ports.
           in_port_base_addr = in_port_base_addr + 'h400;
           if (ingress_ovfl_mode)
              check_probe (.base_addr(in_port_base_addr), .exp_pkt_cnt(exp_ovfl_pkts), .exp_byte_cnt(exp_ovfl_bytes));
           else	   
              check_probe (.base_addr(in_port_base_addr), .exp_pkt_cnt(0), .exp_byte_cnt(0));
        end

        if ( (out_port != HOST_PORT0) ) begin  // no ovfl counters for these egress ports.
           out_port_base_addr = out_port_base_addr + 'h400;
           if (ingress_ovfl_mode)
              check_probe (.base_addr(out_port_base_addr), .exp_pkt_cnt(0), .exp_byte_cnt(0));
           else
              check_probe (.base_addr(out_port_base_addr), .exp_pkt_cnt(exp_ovfl_pkts), .exp_byte_cnt(exp_ovfl_bytes));
        end
       
    endtask;


    task check_err_probes ( input port_t in_port, 
                            input logic [63:0] exp_err_pkts, exp_err_bytes );

        cntr_addr_t in_port_err_addr;
        // establish addr for ingress err counts
        case (in_port)
               CMAC_PORT0 : in_port_err_addr = 'h8800;
               CMAC_PORT1 : in_port_err_addr = 'h9400;
	    default : in_port_err_addr = 'hxxxx;
        endcase

        check_probe (.base_addr(in_port_err_addr), .exp_pkt_cnt(exp_err_pkts), .exp_byte_cnt(exp_err_bytes));

    endtask;


    task check_probe (input cntr_addr_t base_addr, input logic [63:0] exp_pkt_cnt, exp_byte_cnt);
        logic [63:0] rd_data;

        env.reg_agent.read_reg( base_addr + 'h0, rd_data[63:32] );  // pkt_count_upper
        env.reg_agent.read_reg( base_addr + 'h4, rd_data[31:0]  );  // pkt_count_lower
       `INFO($sformatf("%s pkt count: %0d", base_addr.encoded.name(), rd_data));
       `FAIL_UNLESS( rd_data == exp_pkt_cnt );

        env.reg_agent.read_reg( base_addr + 'h8, rd_data[63:32] );  // byte_count_upper
        env.reg_agent.read_reg( base_addr + 'hc, rd_data[31:0]  );  // byte_count_lower
       `INFO($sformatf("%s byte count: %0d", base_addr.encoded.name(), rd_data));
       `FAIL_UNLESS( rd_data == exp_byte_cnt );

    endtask;


    task halt_probe_counters;
        logic [31:0] rd_data;
        bit 	     rd_fail = 0;

        // check initial values.       
        env.probe_from_cmac_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_from_cmac_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_from_host_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_from_host_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);

        env.probe_core_to_app_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_app_to_core_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);

        env.probe_to_cmac_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_to_cmac_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_to_host_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
        env.probe_to_host_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 0);
       `FAIL_UNLESS( rd_fail == 0 );
       
        // set halt_counters.
        env.probe_from_cmac_0_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_from_cmac_1_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_from_host_0_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_from_host_1_reg_blk_agent.write_halt_counters( 8'd1 );

        env.probe_core_to_app_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_app_to_core_reg_blk_agent.write_halt_counters( 8'd1 );

        env.probe_to_cmac_0_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_to_cmac_1_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_to_host_0_reg_blk_agent.write_halt_counters( 8'd1 );
        env.probe_to_host_1_reg_blk_agent.write_halt_counters( 8'd1 );

        // check halt_counters values.
        env.probe_from_cmac_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_from_cmac_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_from_host_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_from_host_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);

        env.probe_core_to_app_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_app_to_core_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);

        env.probe_to_cmac_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_to_cmac_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_to_host_0_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
        env.probe_to_host_1_reg_blk_agent.read_halt_counters( rd_data ); rd_fail = rd_fail || (rd_data != 1);
       `FAIL_UNLESS( rd_fail == 0 );
       
    endtask;
   
endmodule
