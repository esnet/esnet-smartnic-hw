package vitisnetp4_igr_verif_pkg;

   `include "vitisnetp4_igr_agent.svh"

endpackage : vitisnetp4_igr_verif_pkg

