package p4_proc_verif_pkg;
    import p4_proc_reg_verif_pkg::*;

   `include "p4_proc_reg_agent.svh"

endpackage : p4_proc_verif_pkg

