package p4_and_verilog_verif_pkg;
    import p4_and_verilog_reg_verif_pkg::*;

   `include "p4_and_verilog_reg_agent.svh"

endpackage : p4_and_verilog_verif_pkg

