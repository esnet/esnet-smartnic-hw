../../../../../../src/vitisnetp4/verif/include/vitisnetp4_agent.svh