package xilinx_hbm_verif_pkg;

    import xilinx_hbm_reg_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "xilinx_hbm_reg_agent.svh"

endpackage : xilinx_hbm_verif_pkg
