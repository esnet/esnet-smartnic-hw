package xilinx_axis_pkg;

    typedef enum int {
        FULL,
        LITE
    } xilinx_axis_ila_mode_t;

endpackage : xilinx_axis_pkg
