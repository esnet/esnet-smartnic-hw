module xilinx_hbm_stack_if
    import xilinx_hbm_pkg::*;
#(
    parameter density_t DENSITY = DENSITY_4G,
    // Derived parameters (don't override)
    parameter int ADDR_WID = get_addr_wid(DENSITY)
)(
    // Proprietary HBM interface
    // -----------------------------------------
    // HBM reference clock
    input wire logic            hbm_ref_clk,

    // AXI3 memory channel interfaces (16 pseudochannels per stack)
    axi3_intf.peripheral        axi_if [PSEUDO_CHANNELS_PER_STACK],
    
    // APB (management) interface
    apb_intf.peripheral         apb_if,

    // Status
    output wire logic           init_done,
    
    // DRAM status monitoring
    output wire logic           dram_status_cattrip,
    output wire logic [6:0]     dram_status_temp,

    // Xilinx HBM IP (single stack) ports
    // -----------------------------------------
    // Reference clock
    output wire logic                         HBM_REF_CLK_0,
    // Channel 0
    output wire logic                         AXI_00_ACLK,
    output wire logic                         AXI_00_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_00_ARADDR,
    output wire logic [1:0]                   AXI_00_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_00_ARID,
    output wire logic [3:0]                   AXI_00_ARLEN,
    output wire logic [2:0]                   AXI_00_ARSIZE,
    output wire logic                         AXI_00_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_00_AWADDR,
    output wire logic [1:0]                   AXI_00_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_00_AWID,
    output wire logic [3:0]                   AXI_00_AWLEN,
    output wire logic [2:0]                   AXI_00_AWSIZE,
    output wire logic                         AXI_00_AWVALID,
    output wire logic                         AXI_00_RREADY,
    output wire logic                         AXI_00_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_00_WDATA,
    output wire logic                         AXI_00_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_00_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_00_WDATA_PARITY,
    output wire logic                         AXI_00_WVALID,
    input  wire logic                         AXI_00_ARREADY,
    input  wire logic                         AXI_00_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_00_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_00_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_00_RID,
    input  wire logic                         AXI_00_RLAST,
    input  wire logic [1:0]                   AXI_00_RRESP,
    input  wire logic                         AXI_00_RVALID,
    input  wire logic                         AXI_00_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_00_BID,
    input  wire logic [1:0]                   AXI_00_BRESP,
    input  wire logic                         AXI_00_BVALID,
    // Channel 1
    output wire logic                         AXI_01_ACLK,
    output wire logic                         AXI_01_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_01_ARADDR,
    output wire logic [1:0]                   AXI_01_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_01_ARID,
    output wire logic [3:0]                   AXI_01_ARLEN,
    output wire logic [2:0]                   AXI_01_ARSIZE,
    output wire logic                         AXI_01_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_01_AWADDR,
    output wire logic [1:0]                   AXI_01_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_01_AWID,
    output wire logic [3:0]                   AXI_01_AWLEN,
    output wire logic [2:0]                   AXI_01_AWSIZE,
    output wire logic                         AXI_01_AWVALID,
    output wire logic                         AXI_01_RREADY,
    output wire logic                         AXI_01_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_01_WDATA,
    output wire logic                         AXI_01_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_01_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_01_WDATA_PARITY,
    output wire logic                         AXI_01_WVALID,
    input  wire logic                         AXI_01_ARREADY,
    input  wire logic                         AXI_01_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_01_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_01_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_01_RID,
    input  wire logic                         AXI_01_RLAST,
    input  wire logic [1:0]                   AXI_01_RRESP,
    input  wire logic                         AXI_01_RVALID,
    input  wire logic                         AXI_01_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_01_BID,
    input  wire logic [1:0]                   AXI_01_BRESP,
    input  wire logic                         AXI_01_BVALID,
    // Channel 2
    output wire logic                         AXI_02_ACLK,
    output wire logic                         AXI_02_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_02_ARADDR,
    output wire logic [1:0]                   AXI_02_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_02_ARID,
    output wire logic [3:0]                   AXI_02_ARLEN,
    output wire logic [2:0]                   AXI_02_ARSIZE,
    output wire logic                         AXI_02_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_02_AWADDR,
    output wire logic [1:0]                   AXI_02_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_02_AWID,
    output wire logic [3:0]                   AXI_02_AWLEN,
    output wire logic [2:0]                   AXI_02_AWSIZE,
    output wire logic                         AXI_02_AWVALID,
    output wire logic                         AXI_02_RREADY,
    output wire logic                         AXI_02_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_02_WDATA,
    output wire logic                         AXI_02_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_02_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_02_WDATA_PARITY,
    output wire logic                         AXI_02_WVALID,
    input  wire logic                         AXI_02_ARREADY,
    input  wire logic                         AXI_02_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_02_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_02_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_02_RID,
    input  wire logic                         AXI_02_RLAST,
    input  wire logic [1:0]                   AXI_02_RRESP,
    input  wire logic                         AXI_02_RVALID,
    input  wire logic                         AXI_02_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_02_BID,
    input  wire logic [1:0]                   AXI_02_BRESP,
    input  wire logic                         AXI_02_BVALID,
    // Channel 3
    output wire logic                         AXI_03_ACLK,
    output wire logic                         AXI_03_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_03_ARADDR,
    output wire logic [1:0]                   AXI_03_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_03_ARID,
    output wire logic [3:0]                   AXI_03_ARLEN,
    output wire logic [2:0]                   AXI_03_ARSIZE,
    output wire logic                         AXI_03_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_03_AWADDR,
    output wire logic [1:0]                   AXI_03_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_03_AWID,
    output wire logic [3:0]                   AXI_03_AWLEN,
    output wire logic [2:0]                   AXI_03_AWSIZE,
    output wire logic                         AXI_03_AWVALID,
    output wire logic                         AXI_03_RREADY,
    output wire logic                         AXI_03_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_03_WDATA,
    output wire logic                         AXI_03_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_03_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_03_WDATA_PARITY,
    output wire logic                         AXI_03_WVALID,
    input  wire logic                         AXI_03_ARREADY,
    input  wire logic                         AXI_03_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_03_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_03_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_03_RID,
    input  wire logic                         AXI_03_RLAST,
    input  wire logic [1:0]                   AXI_03_RRESP,
    input  wire logic                         AXI_03_RVALID,
    input  wire logic                         AXI_03_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_03_BID,
    input  wire logic [1:0]                   AXI_03_BRESP,
    input  wire logic                         AXI_03_BVALID,
    // Channel 4
    output wire logic                         AXI_04_ACLK,
    output wire logic                         AXI_04_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_04_ARADDR,
    output wire logic [1:0]                   AXI_04_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_04_ARID,
    output wire logic [3:0]                   AXI_04_ARLEN,
    output wire logic [2:0]                   AXI_04_ARSIZE,
    output wire logic                         AXI_04_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_04_AWADDR,
    output wire logic [1:0]                   AXI_04_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_04_AWID,
    output wire logic [3:0]                   AXI_04_AWLEN,
    output wire logic [2:0]                   AXI_04_AWSIZE,
    output wire logic                         AXI_04_AWVALID,
    output wire logic                         AXI_04_RREADY,
    output wire logic                         AXI_04_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_04_WDATA,
    output wire logic                         AXI_04_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_04_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_04_WDATA_PARITY,
    output wire logic                         AXI_04_WVALID,
    input  wire logic                         AXI_04_ARREADY,
    input  wire logic                         AXI_04_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_04_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_04_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_04_RID,
    input  wire logic                         AXI_04_RLAST,
    input  wire logic [1:0]                   AXI_04_RRESP,
    input  wire logic                         AXI_04_RVALID,
    input  wire logic                         AXI_04_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_04_BID,
    input  wire logic [1:0]                   AXI_04_BRESP,
    input  wire logic                         AXI_04_BVALID,
    // Channel 5
    output wire logic                         AXI_05_ACLK,
    output wire logic                         AXI_05_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_05_ARADDR,
    output wire logic [1:0]                   AXI_05_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_05_ARID,
    output wire logic [3:0]                   AXI_05_ARLEN,
    output wire logic [2:0]                   AXI_05_ARSIZE,
    output wire logic                         AXI_05_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_05_AWADDR,
    output wire logic [1:0]                   AXI_05_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_05_AWID,
    output wire logic [3:0]                   AXI_05_AWLEN,
    output wire logic [2:0]                   AXI_05_AWSIZE,
    output wire logic                         AXI_05_AWVALID,
    output wire logic                         AXI_05_RREADY,
    output wire logic                         AXI_05_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_05_WDATA,
    output wire logic                         AXI_05_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_05_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_05_WDATA_PARITY,
    output wire logic                         AXI_05_WVALID,
    input  wire logic                         AXI_05_ARREADY,
    input  wire logic                         AXI_05_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_05_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_05_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_05_RID,
    input  wire logic                         AXI_05_RLAST,
    input  wire logic [1:0]                   AXI_05_RRESP,
    input  wire logic                         AXI_05_RVALID,
    input  wire logic                         AXI_05_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_05_BID,
    input  wire logic [1:0]                   AXI_05_BRESP,
    input  wire logic                         AXI_05_BVALID,
    // Channel 6
    output wire logic                         AXI_06_ACLK,
    output wire logic                         AXI_06_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_06_ARADDR,
    output wire logic [1:0]                   AXI_06_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_06_ARID,
    output wire logic [3:0]                   AXI_06_ARLEN,
    output wire logic [2:0]                   AXI_06_ARSIZE,
    output wire logic                         AXI_06_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_06_AWADDR,
    output wire logic [1:0]                   AXI_06_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_06_AWID,
    output wire logic [3:0]                   AXI_06_AWLEN,
    output wire logic [2:0]                   AXI_06_AWSIZE,
    output wire logic                         AXI_06_AWVALID,
    output wire logic                         AXI_06_RREADY,
    output wire logic                         AXI_06_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_06_WDATA,
    output wire logic                         AXI_06_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_06_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_06_WDATA_PARITY,
    output wire logic                         AXI_06_WVALID,
    input  wire logic                         AXI_06_ARREADY,
    input  wire logic                         AXI_06_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_06_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_06_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_06_RID,
    input  wire logic                         AXI_06_RLAST,
    input  wire logic [1:0]                   AXI_06_RRESP,
    input  wire logic                         AXI_06_RVALID,
    input  wire logic                         AXI_06_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_06_BID,
    input  wire logic [1:0]                   AXI_06_BRESP,
    input  wire logic                         AXI_06_BVALID,
    // Channel 7
    output wire logic                         AXI_07_ACLK,
    output wire logic                         AXI_07_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_07_ARADDR,
    output wire logic [1:0]                   AXI_07_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_07_ARID,
    output wire logic [3:0]                   AXI_07_ARLEN,
    output wire logic [2:0]                   AXI_07_ARSIZE,
    output wire logic                         AXI_07_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_07_AWADDR,
    output wire logic [1:0]                   AXI_07_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_07_AWID,
    output wire logic [3:0]                   AXI_07_AWLEN,
    output wire logic [2:0]                   AXI_07_AWSIZE,
    output wire logic                         AXI_07_AWVALID,
    output wire logic                         AXI_07_RREADY,
    output wire logic                         AXI_07_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_07_WDATA,
    output wire logic                         AXI_07_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_07_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_07_WDATA_PARITY,
    output wire logic                         AXI_07_WVALID,
    input  wire logic                         AXI_07_ARREADY,
    input  wire logic                         AXI_07_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_07_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_07_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_07_RID,
    input  wire logic                         AXI_07_RLAST,
    input  wire logic [1:0]                   AXI_07_RRESP,
    input  wire logic                         AXI_07_RVALID,
    input  wire logic                         AXI_07_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_07_BID,
    input  wire logic [1:0]                   AXI_07_BRESP,
    input  wire logic                         AXI_07_BVALID,
    // Channel 8
    output wire logic                         AXI_08_ACLK,
    output wire logic                         AXI_08_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_08_ARADDR,
    output wire logic [1:0]                   AXI_08_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_08_ARID,
    output wire logic [3:0]                   AXI_08_ARLEN,
    output wire logic [2:0]                   AXI_08_ARSIZE,
    output wire logic                         AXI_08_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_08_AWADDR,
    output wire logic [1:0]                   AXI_08_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_08_AWID,
    output wire logic [3:0]                   AXI_08_AWLEN,
    output wire logic [2:0]                   AXI_08_AWSIZE,
    output wire logic                         AXI_08_AWVALID,
    output wire logic                         AXI_08_RREADY,
    output wire logic                         AXI_08_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_08_WDATA,
    output wire logic                         AXI_08_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_08_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_08_WDATA_PARITY,
    output wire logic                         AXI_08_WVALID,
    input  wire logic                         AXI_08_ARREADY,
    input  wire logic                         AXI_08_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_08_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_08_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_08_RID,
    input  wire logic                         AXI_08_RLAST,
    input  wire logic [1:0]                   AXI_08_RRESP,
    input  wire logic                         AXI_08_RVALID,
    input  wire logic                         AXI_08_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_08_BID,
    input  wire logic [1:0]                   AXI_08_BRESP,
    input  wire logic                         AXI_08_BVALID,
    // Channel 9
    output wire logic                         AXI_09_ACLK,
    output wire logic                         AXI_09_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_09_ARADDR,
    output wire logic [1:0]                   AXI_09_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_09_ARID,
    output wire logic [3:0]                   AXI_09_ARLEN,
    output wire logic [2:0]                   AXI_09_ARSIZE,
    output wire logic                         AXI_09_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_09_AWADDR,
    output wire logic [1:0]                   AXI_09_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_09_AWID,
    output wire logic [3:0]                   AXI_09_AWLEN,
    output wire logic [2:0]                   AXI_09_AWSIZE,
    output wire logic                         AXI_09_AWVALID,
    output wire logic                         AXI_09_RREADY,
    output wire logic                         AXI_09_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_09_WDATA,
    output wire logic                         AXI_09_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_09_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_09_WDATA_PARITY,
    output wire logic                         AXI_09_WVALID,
    input  wire logic                         AXI_09_ARREADY,
    input  wire logic                         AXI_09_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_09_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_09_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_09_RID,
    input  wire logic                         AXI_09_RLAST,
    input  wire logic [1:0]                   AXI_09_RRESP,
    input  wire logic                         AXI_09_RVALID,
    input  wire logic                         AXI_09_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_09_BID,
    input  wire logic [1:0]                   AXI_09_BRESP,
    input  wire logic                         AXI_09_BVALID,
    // Channel 10
    output wire logic                         AXI_10_ACLK,
    output wire logic                         AXI_10_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_10_ARADDR,
    output wire logic [1:0]                   AXI_10_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_10_ARID,
    output wire logic [3:0]                   AXI_10_ARLEN,
    output wire logic [2:0]                   AXI_10_ARSIZE,
    output wire logic                         AXI_10_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_10_AWADDR,
    output wire logic [1:0]                   AXI_10_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_10_AWID,
    output wire logic [3:0]                   AXI_10_AWLEN,
    output wire logic [2:0]                   AXI_10_AWSIZE,
    output wire logic                         AXI_10_AWVALID,
    output wire logic                         AXI_10_RREADY,
    output wire logic                         AXI_10_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_10_WDATA,
    output wire logic                         AXI_10_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_10_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_10_WDATA_PARITY,
    output wire logic                         AXI_10_WVALID,
    input  wire logic                         AXI_10_ARREADY,
    input  wire logic                         AXI_10_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_10_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_10_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_10_RID,
    input  wire logic                         AXI_10_RLAST,
    input  wire logic [1:0]                   AXI_10_RRESP,
    input  wire logic                         AXI_10_RVALID,
    input  wire logic                         AXI_10_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_10_BID,
    input  wire logic [1:0]                   AXI_10_BRESP,
    input  wire logic                         AXI_10_BVALID,
    // Channel 11
    output wire logic                         AXI_11_ACLK,
    output wire logic                         AXI_11_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_11_ARADDR,
    output wire logic [1:0]                   AXI_11_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_11_ARID,
    output wire logic [3:0]                   AXI_11_ARLEN,
    output wire logic [2:0]                   AXI_11_ARSIZE,
    output wire logic                         AXI_11_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_11_AWADDR,
    output wire logic [1:0]                   AXI_11_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_11_AWID,
    output wire logic [3:0]                   AXI_11_AWLEN,
    output wire logic [2:0]                   AXI_11_AWSIZE,
    output wire logic                         AXI_11_AWVALID,
    output wire logic                         AXI_11_RREADY,
    output wire logic                         AXI_11_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_11_WDATA,
    output wire logic                         AXI_11_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_11_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_11_WDATA_PARITY,
    output wire logic                         AXI_11_WVALID,
    input  wire logic                         AXI_11_ARREADY,
    input  wire logic                         AXI_11_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_11_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_11_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_11_RID,
    input  wire logic                         AXI_11_RLAST,
    input  wire logic [1:0]                   AXI_11_RRESP,
    input  wire logic                         AXI_11_RVALID,
    input  wire logic                         AXI_11_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_11_BID,
    input  wire logic [1:0]                   AXI_11_BRESP,
    input  wire logic                         AXI_11_BVALID,
    // Channel 12
    output wire logic                         AXI_12_ACLK,
    output wire logic                         AXI_12_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_12_ARADDR,
    output wire logic [1:0]                   AXI_12_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_12_ARID,
    output wire logic [3:0]                   AXI_12_ARLEN,
    output wire logic [2:0]                   AXI_12_ARSIZE,
    output wire logic                         AXI_12_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_12_AWADDR,
    output wire logic [1:0]                   AXI_12_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_12_AWID,
    output wire logic [3:0]                   AXI_12_AWLEN,
    output wire logic [2:0]                   AXI_12_AWSIZE,
    output wire logic                         AXI_12_AWVALID,
    output wire logic                         AXI_12_RREADY,
    output wire logic                         AXI_12_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_12_WDATA,
    output wire logic                         AXI_12_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_12_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_12_WDATA_PARITY,
    output wire logic                         AXI_12_WVALID,
    input  wire logic                         AXI_12_ARREADY,
    input  wire logic                         AXI_12_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_12_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_12_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_12_RID,
    input  wire logic                         AXI_12_RLAST,
    input  wire logic [1:0]                   AXI_12_RRESP,
    input  wire logic                         AXI_12_RVALID,
    input  wire logic                         AXI_12_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_12_BID,
    input  wire logic [1:0]                   AXI_12_BRESP,
    input  wire logic                         AXI_12_BVALID,
    // Channel 13
    output wire logic                         AXI_13_ACLK,
    output wire logic                         AXI_13_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_13_ARADDR,
    output wire logic [1:0]                   AXI_13_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_13_ARID,
    output wire logic [3:0]                   AXI_13_ARLEN,
    output wire logic [2:0]                   AXI_13_ARSIZE,
    output wire logic                         AXI_13_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_13_AWADDR,
    output wire logic [1:0]                   AXI_13_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_13_AWID,
    output wire logic [3:0]                   AXI_13_AWLEN,
    output wire logic [2:0]                   AXI_13_AWSIZE,
    output wire logic                         AXI_13_AWVALID,
    output wire logic                         AXI_13_RREADY,
    output wire logic                         AXI_13_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_13_WDATA,
    output wire logic                         AXI_13_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_13_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_13_WDATA_PARITY,
    output wire logic                         AXI_13_WVALID,
    input  wire logic                         AXI_13_ARREADY,
    input  wire logic                         AXI_13_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_13_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_13_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_13_RID,
    input  wire logic                         AXI_13_RLAST,
    input  wire logic [1:0]                   AXI_13_RRESP,
    input  wire logic                         AXI_13_RVALID,
    input  wire logic                         AXI_13_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_13_BID,
    input  wire logic [1:0]                   AXI_13_BRESP,
    input  wire logic                         AXI_13_BVALID,
    // Channel 14
    output wire logic                         AXI_14_ACLK,
    output wire logic                         AXI_14_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_14_ARADDR,
    output wire logic [1:0]                   AXI_14_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_14_ARID,
    output wire logic [3:0]                   AXI_14_ARLEN,
    output wire logic [2:0]                   AXI_14_ARSIZE,
    output wire logic                         AXI_14_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_14_AWADDR,
    output wire logic [1:0]                   AXI_14_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_14_AWID,
    output wire logic [3:0]                   AXI_14_AWLEN,
    output wire logic [2:0]                   AXI_14_AWSIZE,
    output wire logic                         AXI_14_AWVALID,
    output wire logic                         AXI_14_RREADY,
    output wire logic                         AXI_14_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_14_WDATA,
    output wire logic                         AXI_14_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_14_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_14_WDATA_PARITY,
    output wire logic                         AXI_14_WVALID,
    input  wire logic                         AXI_14_ARREADY,
    input  wire logic                         AXI_14_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_14_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_14_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_14_RID,
    input  wire logic                         AXI_14_RLAST,
    input  wire logic [1:0]                   AXI_14_RRESP,
    input  wire logic                         AXI_14_RVALID,
    input  wire logic                         AXI_14_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_14_BID,
    input  wire logic [1:0]                   AXI_14_BRESP,
    input  wire logic                         AXI_14_BVALID,
    // Channel 15
    output wire logic                         AXI_15_ACLK,
    output wire logic                         AXI_15_ARESET_N,
    output wire logic [ADDR_WID-1:0]          AXI_15_ARADDR,
    output wire logic [1:0]                   AXI_15_ARBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_15_ARID,
    output wire logic [3:0]                   AXI_15_ARLEN,
    output wire logic [2:0]                   AXI_15_ARSIZE,
    output wire logic                         AXI_15_ARVALID,
    output wire logic [ADDR_WID-1:0]          AXI_15_AWADDR,
    output wire logic [1:0]                   AXI_15_AWBURST,
    output wire logic [AXI_ID_WID-1:0]        AXI_15_AWID,
    output wire logic [3:0]                   AXI_15_AWLEN,
    output wire logic [2:0]                   AXI_15_AWSIZE,
    output wire logic                         AXI_15_AWVALID,
    output wire logic                         AXI_15_RREADY,
    output wire logic                         AXI_15_BREADY,
    output wire logic [AXI_DATA_WID-1:0]      AXI_15_WDATA,
    output wire logic                         AXI_15_WLAST,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_15_WSTRB,
    output wire logic [AXI_DATA_BYTE_WID-1:0] AXI_15_WDATA_PARITY,
    output wire logic                         AXI_15_WVALID,
    input  wire logic                         AXI_15_ARREADY,
    input  wire logic                         AXI_15_AWREADY,
    input  wire logic [AXI_DATA_BYTE_WID-1:0] AXI_15_RDATA_PARITY,
    input  wire logic [AXI_DATA_WID-1:0]      AXI_15_RDATA,
    input  wire logic [AXI_ID_WID-1:0]        AXI_15_RID,
    input  wire logic                         AXI_15_RLAST,
    input  wire logic [1:0]                   AXI_15_RRESP,
    input  wire logic                         AXI_15_RVALID,
    input  wire logic                         AXI_15_WREADY,
    input  wire logic [AXI_ID_WID-1:0]        AXI_15_BID,
    input  wire logic [1:0]                   AXI_15_BRESP,
    input  wire logic                         AXI_15_BVALID,
    // APB interface
    output wire logic [31:0]                  APB_0_PWDATA,
    output wire logic [21:0]                  APB_0_PADDR,
    output wire logic                         APB_0_PCLK,
    output wire logic                         APB_0_PENABLE,
    output wire logic                         APB_0_PRESET_N,
    output wire logic                         APB_0_PSEL,
    output wire logic                         APB_0_PWRITE,
    input  wire logic [31:0]                  APB_0_PRDATA,
    input  wire logic                         APB_0_PREADY,
    input  wire logic                         APB_0_PSLVERR,
    input  wire logic                         apb_complete_0,
    // DRAM status
    input  wire logic                         DRAM_0_STAT_CATTRIP,
    input  wire logic [6:0]                   DRAM_0_STAT_TEMP
);

    // ---------------------------------------
    // Map from wrapper interface to raw IP
    // ---------------------------------------
    // Clock
    assign HBM_REF_CLK_0 = hbm_ref_clk;

    // DRAM status
    assign dram_status_cattrip = DRAM_0_STAT_CATTRIP;
    assign dram_status_temp    = DRAM_0_STAT_TEMP;

    // APB
    apb_intf_to_signals #(
        .DATA_BYTE_WID ( 4 ),
        .ADDR_WID      ( 22 )
    ) i_apb_intf_to_signals (
        .apb_if  ( apb_if ),
        .pclk    ( APB_0_PCLK ),
        .presetn ( APB_0_PRESET_N ),
        .paddr   ( APB_0_PADDR ),
        .pprot   ( ),
        .psel    ( APB_0_PSEL ),
        .penable ( APB_0_PENABLE ),
        .pwrite  ( APB_0_PWRITE ),
        .pwdata  ( APB_0_PWDATA ),
        .pstrb   ( ),
        .pready  ( APB_0_PREADY ),
        .prdata  ( APB_0_PRDATA ),
        .pslverr ( APB_0_PSLVERR )
    );

    assign init_done = apb_complete_0;

    // Memory Channel 0
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch0 (
        .axi3_if  ( axi_if[0] ),
        .aclk     ( AXI_00_ACLK ),
        .aresetn  ( AXI_00_ARESET_N ),
        .awid     ( AXI_00_AWID ),
        .awaddr   ( AXI_00_AWADDR ),
        .awlen    ( AXI_00_AWLEN ),
        .awsize   ( AXI_00_AWSIZE ),
        .awburst  ( AXI_00_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_00_AWVALID ),
        .awready  ( AXI_00_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_00_WDATA ),
        .wstrb    ( AXI_00_WSTRB ),
        .wlast    ( AXI_00_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_00_WVALID ),
        .wready   ( AXI_00_WREADY ),
        .bid      ( AXI_00_BID ),
        .bresp    ( AXI_00_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_00_BVALID ),
        .bready   ( AXI_00_BREADY ),
        .arid     ( AXI_00_ARID ),
        .araddr   ( AXI_00_ARADDR ),
        .arlen    ( AXI_00_ARLEN ),
        .arsize   ( AXI_00_ARSIZE ),
        .arburst  ( AXI_00_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_00_ARVALID ),
        .arready  ( AXI_00_ARREADY ),
        .rid      ( AXI_00_RID ),
        .rdata    ( AXI_00_RDATA ),
        .rresp    ( AXI_00_RRESP ),
        .rlast    ( AXI_00_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_00_RVALID ),
        .rready   ( AXI_00_RREADY )
    );

    assign AXI_00_WDATA_PARITY = '0;
  
    // Memory Channel 1
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch1 (
        .axi3_if  ( axi_if[1] ),
        .aclk     ( AXI_01_ACLK ),
        .aresetn  ( AXI_01_ARESET_N ),
        .awid     ( AXI_01_AWID ),
        .awaddr   ( AXI_01_AWADDR ),
        .awlen    ( AXI_01_AWLEN ),
        .awsize   ( AXI_01_AWSIZE ),
        .awburst  ( AXI_01_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_01_AWVALID ),
        .awready  ( AXI_01_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_01_WDATA ),
        .wstrb    ( AXI_01_WSTRB ),
        .wlast    ( AXI_01_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_01_WVALID ),
        .wready   ( AXI_01_WREADY ),
        .bid      ( AXI_01_BID ),
        .bresp    ( AXI_01_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_01_BVALID ),
        .bready   ( AXI_01_BREADY ),
        .arid     ( AXI_01_ARID ),
        .araddr   ( AXI_01_ARADDR ),
        .arlen    ( AXI_01_ARLEN ),
        .arsize   ( AXI_01_ARSIZE ),
        .arburst  ( AXI_01_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_01_ARVALID ),
        .arready  ( AXI_01_ARREADY ),
        .rid      ( AXI_01_RID ),
        .rdata    ( AXI_01_RDATA ),
        .rresp    ( AXI_01_RRESP ),
        .rlast    ( AXI_01_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_01_RVALID ),
        .rready   ( AXI_01_RREADY )
    );

    assign AXI_01_WDATA_PARITY = '0;
 
    // Memory Channel 2
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch2 (
        .axi3_if  ( axi_if[2] ),
        .aclk     ( AXI_02_ACLK ),
        .aresetn  ( AXI_02_ARESET_N ),
        .awid     ( AXI_02_AWID ),
        .awaddr   ( AXI_02_AWADDR ),
        .awlen    ( AXI_02_AWLEN ),
        .awsize   ( AXI_02_AWSIZE ),
        .awburst  ( AXI_02_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_02_AWVALID ),
        .awready  ( AXI_02_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_02_WDATA ),
        .wstrb    ( AXI_02_WSTRB ),
        .wlast    ( AXI_02_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_02_WVALID ),
        .wready   ( AXI_02_WREADY ),
        .bid      ( AXI_02_BID ),
        .bresp    ( AXI_02_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_02_BVALID ),
        .bready   ( AXI_02_BREADY ),
        .arid     ( AXI_02_ARID ),
        .araddr   ( AXI_02_ARADDR ),
        .arlen    ( AXI_02_ARLEN ),
        .arsize   ( AXI_02_ARSIZE ),
        .arburst  ( AXI_02_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_02_ARVALID ),
        .arready  ( AXI_02_ARREADY ),
        .rid      ( AXI_02_RID ),
        .rdata    ( AXI_02_RDATA ),
        .rresp    ( AXI_02_RRESP ),
        .rlast    ( AXI_02_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_02_RVALID ),
        .rready   ( AXI_02_RREADY )
    );

    assign AXI_02_WDATA_PARITY = '0;
 
    // Memory Channel 3
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch3 (
        .axi3_if  ( axi_if[3] ),
        .aclk     ( AXI_03_ACLK ),
        .aresetn  ( AXI_03_ARESET_N ),
        .awid     ( AXI_03_AWID ),
        .awaddr   ( AXI_03_AWADDR ),
        .awlen    ( AXI_03_AWLEN ),
        .awsize   ( AXI_03_AWSIZE ),
        .awburst  ( AXI_03_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_03_AWVALID ),
        .awready  ( AXI_03_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_03_WDATA ),
        .wstrb    ( AXI_03_WSTRB ),
        .wlast    ( AXI_03_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_03_WVALID ),
        .wready   ( AXI_03_WREADY ),
        .bid      ( AXI_03_BID ),
        .bresp    ( AXI_03_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_03_BVALID ),
        .bready   ( AXI_03_BREADY ),
        .arid     ( AXI_03_ARID ),
        .araddr   ( AXI_03_ARADDR ),
        .arlen    ( AXI_03_ARLEN ),
        .arsize   ( AXI_03_ARSIZE ),
        .arburst  ( AXI_03_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_03_ARVALID ),
        .arready  ( AXI_03_ARREADY ),
        .rid      ( AXI_03_RID ),
        .rdata    ( AXI_03_RDATA ),
        .rresp    ( AXI_03_RRESP ),
        .rlast    ( AXI_03_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_03_RVALID ),
        .rready   ( AXI_03_RREADY )
    );

    assign AXI_03_WDATA_PARITY = '0;

    // Memory Channel 4
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch4 (
        .axi3_if  ( axi_if[4] ),
        .aclk     ( AXI_04_ACLK ),
        .aresetn  ( AXI_04_ARESET_N ),
        .awid     ( AXI_04_AWID ),
        .awaddr   ( AXI_04_AWADDR ),
        .awlen    ( AXI_04_AWLEN ),
        .awsize   ( AXI_04_AWSIZE ),
        .awburst  ( AXI_04_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_04_AWVALID ),
        .awready  ( AXI_04_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_04_WDATA ),
        .wstrb    ( AXI_04_WSTRB ),
        .wlast    ( AXI_04_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_04_WVALID ),
        .wready   ( AXI_04_WREADY ),
        .bid      ( AXI_04_BID ),
        .bresp    ( AXI_04_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_04_BVALID ),
        .bready   ( AXI_04_BREADY ),
        .arid     ( AXI_04_ARID ),
        .araddr   ( AXI_04_ARADDR ),
        .arlen    ( AXI_04_ARLEN ),
        .arsize   ( AXI_04_ARSIZE ),
        .arburst  ( AXI_04_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_04_ARVALID ),
        .arready  ( AXI_04_ARREADY ),
        .rid      ( AXI_04_RID ),
        .rdata    ( AXI_04_RDATA ),
        .rresp    ( AXI_04_RRESP ),
        .rlast    ( AXI_04_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_04_RVALID ),
        .rready   ( AXI_04_RREADY )
    );

    assign AXI_04_WDATA_PARITY = '0;
 
    // Memory Channel 5
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch5 (
        .axi3_if  ( axi_if[5] ),
        .aclk     ( AXI_05_ACLK ),
        .aresetn  ( AXI_05_ARESET_N ),
        .awid     ( AXI_05_AWID ),
        .awaddr   ( AXI_05_AWADDR ),
        .awlen    ( AXI_05_AWLEN ),
        .awsize   ( AXI_05_AWSIZE ),
        .awburst  ( AXI_05_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_05_AWVALID ),
        .awready  ( AXI_05_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_05_WDATA ),
        .wstrb    ( AXI_05_WSTRB ),
        .wlast    ( AXI_05_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_05_WVALID ),
        .wready   ( AXI_05_WREADY ),
        .bid      ( AXI_05_BID ),
        .bresp    ( AXI_05_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_05_BVALID ),
        .bready   ( AXI_05_BREADY ),
        .arid     ( AXI_05_ARID ),
        .araddr   ( AXI_05_ARADDR ),
        .arlen    ( AXI_05_ARLEN ),
        .arsize   ( AXI_05_ARSIZE ),
        .arburst  ( AXI_05_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_05_ARVALID ),
        .arready  ( AXI_05_ARREADY ),
        .rid      ( AXI_05_RID ),
        .rdata    ( AXI_05_RDATA ),
        .rresp    ( AXI_05_RRESP ),
        .rlast    ( AXI_05_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_05_RVALID ),
        .rready   ( AXI_05_RREADY )
    );

    assign AXI_05_WDATA_PARITY = '0;

    // Memory Channel 6
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch6 (
        .axi3_if  ( axi_if[6] ),
        .aclk     ( AXI_06_ACLK ),
        .aresetn  ( AXI_06_ARESET_N ),
        .awid     ( AXI_06_AWID ),
        .awaddr   ( AXI_06_AWADDR ),
        .awlen    ( AXI_06_AWLEN ),
        .awsize   ( AXI_06_AWSIZE ),
        .awburst  ( AXI_06_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_06_AWVALID ),
        .awready  ( AXI_06_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_06_WDATA ),
        .wstrb    ( AXI_06_WSTRB ),
        .wlast    ( AXI_06_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_06_WVALID ),
        .wready   ( AXI_06_WREADY ),
        .bid      ( AXI_06_BID ),
        .bresp    ( AXI_06_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_06_BVALID ),
        .bready   ( AXI_06_BREADY ),
        .arid     ( AXI_06_ARID ),
        .araddr   ( AXI_06_ARADDR ),
        .arlen    ( AXI_06_ARLEN ),
        .arsize   ( AXI_06_ARSIZE ),
        .arburst  ( AXI_06_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_06_ARVALID ),
        .arready  ( AXI_06_ARREADY ),
        .rid      ( AXI_06_RID ),
        .rdata    ( AXI_06_RDATA ),
        .rresp    ( AXI_06_RRESP ),
        .rlast    ( AXI_06_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_06_RVALID ),
        .rready   ( AXI_06_RREADY )
    );

    assign AXI_06_WDATA_PARITY = '0;
 
    // Memory Channel 7
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch7 (
        .axi3_if  ( axi_if[7] ),
        .aclk     ( AXI_07_ACLK ),
        .aresetn  ( AXI_07_ARESET_N ),
        .awid     ( AXI_07_AWID ),
        .awaddr   ( AXI_07_AWADDR ),
        .awlen    ( AXI_07_AWLEN ),
        .awsize   ( AXI_07_AWSIZE ),
        .awburst  ( AXI_07_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_07_AWVALID ),
        .awready  ( AXI_07_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_07_WDATA ),
        .wstrb    ( AXI_07_WSTRB ),
        .wlast    ( AXI_07_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_07_WVALID ),
        .wready   ( AXI_07_WREADY ),
        .bid      ( AXI_07_BID ),
        .bresp    ( AXI_07_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_07_BVALID ),
        .bready   ( AXI_07_BREADY ),
        .arid     ( AXI_07_ARID ),
        .araddr   ( AXI_07_ARADDR ),
        .arlen    ( AXI_07_ARLEN ),
        .arsize   ( AXI_07_ARSIZE ),
        .arburst  ( AXI_07_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_07_ARVALID ),
        .arready  ( AXI_07_ARREADY ),
        .rid      ( AXI_07_RID ),
        .rdata    ( AXI_07_RDATA ),
        .rresp    ( AXI_07_RRESP ),
        .rlast    ( AXI_07_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_07_RVALID ),
        .rready   ( AXI_07_RREADY )
    );

    assign AXI_07_WDATA_PARITY = '0;
 
    // Memory Channel 8
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch8 (
        .axi3_if  ( axi_if[8] ),
        .aclk     ( AXI_08_ACLK ),
        .aresetn  ( AXI_08_ARESET_N ),
        .awid     ( AXI_08_AWID ),
        .awaddr   ( AXI_08_AWADDR ),
        .awlen    ( AXI_08_AWLEN ),
        .awsize   ( AXI_08_AWSIZE ),
        .awburst  ( AXI_08_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_08_AWVALID ),
        .awready  ( AXI_08_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_08_WDATA ),
        .wstrb    ( AXI_08_WSTRB ),
        .wlast    ( AXI_08_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_08_WVALID ),
        .wready   ( AXI_08_WREADY ),
        .bid      ( AXI_08_BID ),
        .bresp    ( AXI_08_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_08_BVALID ),
        .bready   ( AXI_08_BREADY ),
        .arid     ( AXI_08_ARID ),
        .araddr   ( AXI_08_ARADDR ),
        .arlen    ( AXI_08_ARLEN ),
        .arsize   ( AXI_08_ARSIZE ),
        .arburst  ( AXI_08_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_08_ARVALID ),
        .arready  ( AXI_08_ARREADY ),
        .rid      ( AXI_08_RID ),
        .rdata    ( AXI_08_RDATA ),
        .rresp    ( AXI_08_RRESP ),
        .rlast    ( AXI_08_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_08_RVALID ),
        .rready   ( AXI_08_RREADY )
    );

    assign AXI_08_WDATA_PARITY = '0;
 
    // Memory Channel 9
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch9 (
        .axi3_if  ( axi_if[9] ),
        .aclk     ( AXI_09_ACLK ),
        .aresetn  ( AXI_09_ARESET_N ),
        .awid     ( AXI_09_AWID ),
        .awaddr   ( AXI_09_AWADDR ),
        .awlen    ( AXI_09_AWLEN ),
        .awsize   ( AXI_09_AWSIZE ),
        .awburst  ( AXI_09_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_09_AWVALID ),
        .awready  ( AXI_09_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_09_WDATA ),
        .wstrb    ( AXI_09_WSTRB ),
        .wlast    ( AXI_09_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_09_WVALID ),
        .wready   ( AXI_09_WREADY ),
        .bid      ( AXI_09_BID ),
        .bresp    ( AXI_09_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_09_BVALID ),
        .bready   ( AXI_09_BREADY ),
        .arid     ( AXI_09_ARID ),
        .araddr   ( AXI_09_ARADDR ),
        .arlen    ( AXI_09_ARLEN ),
        .arsize   ( AXI_09_ARSIZE ),
        .arburst  ( AXI_09_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_09_ARVALID ),
        .arready  ( AXI_09_ARREADY ),
        .rid      ( AXI_09_RID ),
        .rdata    ( AXI_09_RDATA ),
        .rresp    ( AXI_09_RRESP ),
        .rlast    ( AXI_09_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_09_RVALID ),
        .rready   ( AXI_09_RREADY )
    );

    assign AXI_09_WDATA_PARITY = '0;

    // Memory Channel 10
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch10 (
        .axi3_if  ( axi_if[10] ),
        .aclk     ( AXI_10_ACLK ),
        .aresetn  ( AXI_10_ARESET_N ),
        .awid     ( AXI_10_AWID ),
        .awaddr   ( AXI_10_AWADDR ),
        .awlen    ( AXI_10_AWLEN ),
        .awsize   ( AXI_10_AWSIZE ),
        .awburst  ( AXI_10_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_10_AWVALID ),
        .awready  ( AXI_10_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_10_WDATA ),
        .wstrb    ( AXI_10_WSTRB ),
        .wlast    ( AXI_10_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_10_WVALID ),
        .wready   ( AXI_10_WREADY ),
        .bid      ( AXI_10_BID ),
        .bresp    ( AXI_10_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_10_BVALID ),
        .bready   ( AXI_10_BREADY ),
        .arid     ( AXI_10_ARID ),
        .araddr   ( AXI_10_ARADDR ),
        .arlen    ( AXI_10_ARLEN ),
        .arsize   ( AXI_10_ARSIZE ),
        .arburst  ( AXI_10_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_10_ARVALID ),
        .arready  ( AXI_10_ARREADY ),
        .rid      ( AXI_10_RID ),
        .rdata    ( AXI_10_RDATA ),
        .rresp    ( AXI_10_RRESP ),
        .rlast    ( AXI_10_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_10_RVALID ),
        .rready   ( AXI_10_RREADY )
    );

    assign AXI_10_WDATA_PARITY = '0;

    // Memory Channel 11
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch11 (
        .axi3_if  ( axi_if[11] ),
        .aclk     ( AXI_11_ACLK ),
        .aresetn  ( AXI_11_ARESET_N ),
        .awid     ( AXI_11_AWID ),
        .awaddr   ( AXI_11_AWADDR ),
        .awlen    ( AXI_11_AWLEN ),
        .awsize   ( AXI_11_AWSIZE ),
        .awburst  ( AXI_11_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_11_AWVALID ),
        .awready  ( AXI_11_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_11_WDATA ),
        .wstrb    ( AXI_11_WSTRB ),
        .wlast    ( AXI_11_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_11_WVALID ),
        .wready   ( AXI_11_WREADY ),
        .bid      ( AXI_11_BID ),
        .bresp    ( AXI_11_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_11_BVALID ),
        .bready   ( AXI_11_BREADY ),
        .arid     ( AXI_11_ARID ),
        .araddr   ( AXI_11_ARADDR ),
        .arlen    ( AXI_11_ARLEN ),
        .arsize   ( AXI_11_ARSIZE ),
        .arburst  ( AXI_11_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_11_ARVALID ),
        .arready  ( AXI_11_ARREADY ),
        .rid      ( AXI_11_RID ),
        .rdata    ( AXI_11_RDATA ),
        .rresp    ( AXI_11_RRESP ),
        .rlast    ( AXI_11_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_11_RVALID ),
        .rready   ( AXI_11_RREADY )
    );

    assign AXI_11_WDATA_PARITY = '0;

    // Memory Channel 12
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch12 (
        .axi3_if  ( axi_if[12] ),
        .aclk     ( AXI_12_ACLK ),
        .aresetn  ( AXI_12_ARESET_N ),
        .awid     ( AXI_12_AWID ),
        .awaddr   ( AXI_12_AWADDR ),
        .awlen    ( AXI_12_AWLEN ),
        .awsize   ( AXI_12_AWSIZE ),
        .awburst  ( AXI_12_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_12_AWVALID ),
        .awready  ( AXI_12_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_12_WDATA ),
        .wstrb    ( AXI_12_WSTRB ),
        .wlast    ( AXI_12_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_12_WVALID ),
        .wready   ( AXI_12_WREADY ),
        .bid      ( AXI_12_BID ),
        .bresp    ( AXI_12_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_12_BVALID ),
        .bready   ( AXI_12_BREADY ),
        .arid     ( AXI_12_ARID ),
        .araddr   ( AXI_12_ARADDR ),
        .arlen    ( AXI_12_ARLEN ),
        .arsize   ( AXI_12_ARSIZE ),
        .arburst  ( AXI_12_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_12_ARVALID ),
        .arready  ( AXI_12_ARREADY ),
        .rid      ( AXI_12_RID ),
        .rdata    ( AXI_12_RDATA ),
        .rresp    ( AXI_12_RRESP ),
        .rlast    ( AXI_12_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_12_RVALID ),
        .rready   ( AXI_12_RREADY )
    );

    assign AXI_12_WDATA_PARITY = '0;

    // Memory Channel 13
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch13 (
        .axi3_if  ( axi_if[13] ),
        .aclk     ( AXI_13_ACLK ),
        .aresetn  ( AXI_13_ARESET_N ),
        .awid     ( AXI_13_AWID ),
        .awaddr   ( AXI_13_AWADDR ),
        .awlen    ( AXI_13_AWLEN ),
        .awsize   ( AXI_13_AWSIZE ),
        .awburst  ( AXI_13_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_13_AWVALID ),
        .awready  ( AXI_13_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_13_WDATA ),
        .wstrb    ( AXI_13_WSTRB ),
        .wlast    ( AXI_13_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_13_WVALID ),
        .wready   ( AXI_13_WREADY ),
        .bid      ( AXI_13_BID ),
        .bresp    ( AXI_13_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_13_BVALID ),
        .bready   ( AXI_13_BREADY ),
        .arid     ( AXI_13_ARID ),
        .araddr   ( AXI_13_ARADDR ),
        .arlen    ( AXI_13_ARLEN ),
        .arsize   ( AXI_13_ARSIZE ),
        .arburst  ( AXI_13_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_13_ARVALID ),
        .arready  ( AXI_13_ARREADY ),
        .rid      ( AXI_13_RID ),
        .rdata    ( AXI_13_RDATA ),
        .rresp    ( AXI_13_RRESP ),
        .rlast    ( AXI_13_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_13_RVALID ),
        .rready   ( AXI_13_RREADY )
    );

    assign AXI_13_WDATA_PARITY = '0;

    // Memory Channel 14
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch14 (
        .axi3_if  ( axi_if[14] ),
        .aclk     ( AXI_14_ACLK ),
        .aresetn  ( AXI_14_ARESET_N ),
        .awid     ( AXI_14_AWID ),
        .awaddr   ( AXI_14_AWADDR ),
        .awlen    ( AXI_14_AWLEN ),
        .awsize   ( AXI_14_AWSIZE ),
        .awburst  ( AXI_14_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_14_AWVALID ),
        .awready  ( AXI_14_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_14_WDATA ),
        .wstrb    ( AXI_14_WSTRB ),
        .wlast    ( AXI_14_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_14_WVALID ),
        .wready   ( AXI_14_WREADY ),
        .bid      ( AXI_14_BID ),
        .bresp    ( AXI_14_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_14_BVALID ),
        .bready   ( AXI_14_BREADY ),
        .arid     ( AXI_14_ARID ),
        .araddr   ( AXI_14_ARADDR ),
        .arlen    ( AXI_14_ARLEN ),
        .arsize   ( AXI_14_ARSIZE ),
        .arburst  ( AXI_14_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_14_ARVALID ),
        .arready  ( AXI_14_ARREADY ),
        .rid      ( AXI_14_RID ),
        .rdata    ( AXI_14_RDATA ),
        .rresp    ( AXI_14_RRESP ),
        .rlast    ( AXI_14_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_14_RVALID ),
        .rready   ( AXI_14_RREADY )
    );

    assign AXI_14_WDATA_PARITY = '0;

    // Memory Channel 15
    axi3_intf_to_signals #(
        .DATA_BYTE_WID ( 32 ),
        .ADDR_WID      ( ADDR_WID ),
        .ID_WID        ( AXI_ID_WID )
    ) i_axi3_intf_to_signals__ch15 (
        .axi3_if  ( axi_if[15] ),
        .aclk     ( AXI_15_ACLK ),
        .aresetn  ( AXI_15_ARESET_N ),
        .awid     ( AXI_15_AWID ),
        .awaddr   ( AXI_15_AWADDR ),
        .awlen    ( AXI_15_AWLEN ),
        .awsize   ( AXI_15_AWSIZE ),
        .awburst  ( AXI_15_AWBURST ),
        .awlock   ( ),
        .awcache  ( ),
        .awprot   ( ),
        .awqos    ( ),
        .awregion ( ),
        .awuser   ( ),
        .awvalid  ( AXI_15_AWVALID ),
        .awready  ( AXI_15_AWREADY ),
        .wid      ( ),
        .wdata    ( AXI_15_WDATA ),
        .wstrb    ( AXI_15_WSTRB ),
        .wlast    ( AXI_15_WLAST ),
        .wuser    ( ),
        .wvalid   ( AXI_15_WVALID ),
        .wready   ( AXI_15_WREADY ),
        .bid      ( AXI_15_BID ),
        .bresp    ( AXI_15_BRESP ),
        .buser    ( '0 ),
        .bvalid   ( AXI_15_BVALID ),
        .bready   ( AXI_15_BREADY ),
        .arid     ( AXI_15_ARID ),
        .araddr   ( AXI_15_ARADDR ),
        .arlen    ( AXI_15_ARLEN ),
        .arsize   ( AXI_15_ARSIZE ),
        .arburst  ( AXI_15_ARBURST ),
        .arlock   ( ),
        .arcache  ( ),
        .arprot   ( ),
        .arqos    ( ),
        .arregion ( ),
        .aruser   ( ),
        .arvalid  ( AXI_15_ARVALID ),
        .arready  ( AXI_15_ARREADY ),
        .rid      ( AXI_15_RID ),
        .rdata    ( AXI_15_RDATA ),
        .rresp    ( AXI_15_RRESP ),
        .rlast    ( AXI_15_RLAST ),
        .ruser    ( '0 ),
        .rvalid   ( AXI_15_RVALID ),
        .rready   ( AXI_15_RREADY )
    );

    assign AXI_15_WDATA_PARITY = '0;

endmodule : xilinx_hbm_stack_if
