package vitisnetp4_egr_verif_pkg;

   `include "vitisnetp4_egr_agent.svh"

endpackage : vitisnetp4_egr_verif_pkg

