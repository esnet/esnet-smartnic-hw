package smartnic_app_verif_pkg;
    import smartnic_app_p4_only_reg_verif_pkg::*;

   `include "p4_only_reg_agent.svh"

endpackage : smartnic_app_verif_pkg
