package proxy_test_verif_pkg;
    import proxy_test_reg_verif_pkg::*;

   `include "proxy_test_reg_agent.svh"

endpackage : proxy_test_verif_pkg

