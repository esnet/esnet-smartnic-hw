// Application core (black-box version)
// (used for OOC synthesis of shell)
(* black_box *) module core #() (
    // Shell interface
    shell_intf.core shell_if
);
endmodule : core
