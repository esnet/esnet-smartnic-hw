package smartnic_app_verif_pkg;
    import smartnic_app_reg_verif_pkg::*;

   `include "smartnic_app_reg_agent.svh"

endpackage : smartnic_app_verif_pkg
