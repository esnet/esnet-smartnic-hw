package tb_pkg;
    import axi4l_verif_pkg::*;
    import axi4s_verif_pkg::*;
    import smartnic_reg_verif_pkg::*;
    import axi4s_reg_verif_pkg::*;
    import reg_endian_reg_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "tb_env.svh"

endpackage : tb_pkg
