package xilinx_cms_pkg;

endpackage : xilinx_cms_pkg
