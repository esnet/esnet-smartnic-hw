package `VITISNETP4_VERIF_PKG_NAME;

   `include "vitisnetp4_agent.svh"

endpackage : `VITISNETP4_VERIF_PKG_NAME

