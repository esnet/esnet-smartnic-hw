    // AXI4 interface (signals)
    input         axi_clk;
    input         axi_resetn;
    input  [41:0] APP_AXI_araddr;
    input  [1:0]  APP_AXI_arburst;
    input  [3:0]  APP_AXI_arcache;
    input  [7:0]  APP_AXI_arlen;
    input  [0:0]  APP_AXI_arlock;
    input  [2:0]  APP_AXI_arprot;
    input  [3:0]  APP_AXI_arqos;
    output        APP_AXI_arready;
    input  [2:0]  APP_AXI_arsize;
    input  [17:0] APP_AXI_aruser;
    input         APP_AXI_arvalid;
    input  [41:0] APP_AXI_awaddr;
    input  [1:0]  APP_AXI_awburst;
    input  [3:0]  APP_AXI_awcache;
    input  [7:0]  APP_AXI_awlen;
    input  [0:0]  APP_AXI_awlock;
    input  [2:0]  APP_AXI_awprot;
    input  [3:0]  APP_AXI_awqos;
    output        APP_AXI_awready;
    input  [2:0]  APP_AXI_awsize;
    input  [17:0] APP_AXI_awuser;
    input         APP_AXI_awvalid;
    input         APP_AXI_bready;
    output [1:0]  APP_AXI_bresp;
    output        APP_AXI_bvalid;
    output [31:0] APP_AXI_rdata;
    output        APP_AXI_rlast;
    input         APP_AXI_rready;
    output [1:0]  APP_AXI_rresp;
    output        APP_AXI_rvalid;
    input  [31:0] APP_AXI_wdata;
    input         APP_AXI_wlast;
    output        APP_AXI_wready;
    input  [3:0]  APP_AXI_wstrb;
    input         APP_AXI_wvalid;
