package p4_app_verif_pkg;
    import p4_app_reg_verif_pkg::*;

   `include "p4_app_reg_agent.svh"

endpackage : p4_app_verif_pkg

