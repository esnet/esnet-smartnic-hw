// Nothing to do
// - this file is expected by the OpenNIC Shell build script;
//   in the SmartNIC context, the register map is defined
//   in regio so the file is required but the contents are not
