package xilinx_sysmon_pkg;

endpackage : xilinx_sysmon_pkg
