config xilinx_qdma_sim_cfg;
    design xilinx__qdma__rtl.xilinx_qdma_wrapper;
    default liblist unifast_ver;
endconfig
