module smartnic_app_igr_p4_default ();
    // Dummy module to force compilation library creation.
endmodule
