package xilinx_alveo_au55c_pkg;

    // --------------------------------------------------------------
    // Parameters
    // --------------------------------------------------------------
    localparam int PCIE_LINK_WID = 16;
    localparam int NUM_CMAC = 2;

endpackage : xilinx_alveo_au55c_pkg
