package vitisnetp4_verif_pkg;

   `include "vitisnetp4_agent.svh"

endpackage : vitisnetp4_verif_pkg

