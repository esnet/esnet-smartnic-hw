package sdnet_igr_app_pkg;

    localparam bit INCLUDE_HBM = 1'b0;

endpackage : sdnet_igr_app_pkg
