package smartnic_verif_pkg;
    import std_verif_pkg::*;
    import axi4s_verif_pkg::*;
    import reg_endian_reg_verif_pkg::*;
    import smartnic_pkg::*;

    // Testbench class definitions
    // (declared here to enforce smartnic_verif_pkg::* namespace)
    `include "smartnic_model.svh"
    `include "smartnic_env.svh"

endpackage : smartnic_verif_pkg
